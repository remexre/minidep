grammar edu:umn:cs:melt:minidep:util;

function builtin
Location ::=
{
  return txtLoc("builtin");
}
