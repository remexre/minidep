grammar edu:umn:cs:melt:minidep:abstractsyntax:spined;
